library IEEE;
use IEEE.std_logic_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY test3 IS 
END test3;

ARCHITECTURE test OF test3 IS
COMPONENT mult IS
GENERIC(n : INTEGER := 4 );
PORT   (a : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	b : IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
	ANS : OUT STD_LOGIC_VECTOR(2*n - 1 DOWNTO 0));
END COMPONENT;

--FOR ALL: m1 USE ENTITY WORK.mult(BEHAVIORAL);

CONSTANT n4 : INTEGER := 4;
CONSTANT n8 : INTEGER := 8;

SIGNAL x4 , y4: STD_LOGIC_VECTOR(n4-1 DOWNTO 0);
SIGNAL x8 , y8: STD_LOGIC_VECTOR(n8-1 DOWNTO 0);
SIGNAL ans4 : STD_LOGIC_VECTOR(2*n4-1 DOWNTO 0);
SIGNAL ans8 : STD_LOGIC_VECTOR(2*n8-1 DOWNTO 0);

BEGIN 
	TST4 : mult GENERIC MAP(n => n4)
		  PORT MAP(a => x4 , b => y4 , ANS => ans4);
	x4 <= "1101" , "1111" AFTER 100 NS;
	y4 <= "1010" , "1111" AFTER 100 NS;

	TST8 : mult GENERIC MAP(n => n8)
		  PORT MAP(a => x8 , b => y8 , ANS => ans8);
	x8 <= "10000001";
	y8 <= "10101000";
END test;
